module task_test(
    Clk,
    Reset_n,
    a
);
    input Clk;
    input Reset_n;
    input [3:0]a;
endmodule