module DDS_Module_AD9767(
	Clk,
);

endmodule